        // @subst[`echo $SUBST_TEST_ENV_VAR`]
        // @endsubst
