        // @subst[`echo $SUBST_TEST_ENV_VAR`]
        42
        // @endsubst
