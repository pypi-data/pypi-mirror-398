        // @subst[`printf`]
        // @endsubst
