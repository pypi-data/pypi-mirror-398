`ifndef __MULTI_VAR_TEMPLATE_SVH__
`define __MULTI_VAR_TEMPLATE_SVH__

`define PRIMARY_IMAGE_PATH    `"/primary/path/primary_image.hex`"
`define SECONDARY_IMAGE_PATH  `"/secondary/path/secondary_image.hex`"

`endif // __MULTI_VAR_TEMPLATE_SVH__

