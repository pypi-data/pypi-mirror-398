        // @subst[`printf`]
        Hello, world!
        // @endsubst
