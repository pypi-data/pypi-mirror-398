// @subst[`printf "%s\n%d\n" 'hello, world' 999`]
// @endsubst
// @subst[`printf '%d\n%d\n' 888 777`]
// @endsubst