`ifndef __FLASH_DEFINES_SVH__
`define __FLASH_DEFINES_SVH__

`define QSPIFLASH_PAGE_WRITE_BUFFER_HEX    `"/a/b/c/qspiflash_initial_page_buffer_ram.hex`"
`define QSPIFLASHWB_PAGE_WRITE_BUFFER_HEX  `"/a/b/c/qspiflashwb_initial_page_buffer_ram.hex`"
`define QSPIFLASHWB_READ_CACHE_HEX         `"/a/b/c/qspiflashwb_initial_read_cache_ram.hex`"

`endif // __FLASH_DEFINES_SVH__